** sch_path: /home/amedcalf/projects/flash_circuits/sonos/sonos_curves_simple.sch
**.subckt sonos_curves_simple
XM1 vd vg vs vb sky130_fd_bs_flash__special_sonosfet_star L=0.22 W=0.45 nf=1 ad='1 * W * 0.29' as='1 * W * 0.29' pd='2 * (W + 0.29)'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vd vg vs vb sky130_fd_bs_flash__special_sonosfet_original L=0.22 W=0.45 nf=1 ad='1 * W * 0.29' as='1 * W * 0.29' pd='2 * (W + 0.29)'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
vg vg GND 0
vd vd GND 1
vs vs GND 0
vb vb GND 0
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
.include /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sonos_see_e/begin_of_life.spice
.include /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sonos_see_e/begin_of_life.pm3.spice
.include /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sonos_see_p/begin_of_life.spice
.include /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sonos_see_p/begin_of_life.pm3.spice



.option savecurrents
*.option abstol=1e-10 reltol=1e-2 chgtol=1e-12
*.ic v(bootp)=0 v(bootn)=0 v(inp)=0 v(inn)=0 v(inf)=0 v(inb)=0
*.ic v(net3)=0 v(net4)=0
.control
  unset appendwrite
  save all

  dc vd 0 1 0.1 vg 0 2 0.5
  remzerovec
  write test_sonos_curves_simple.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
