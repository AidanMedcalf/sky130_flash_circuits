** sch_path: /home/amedcalf/projects/flash_circuits/row_drivers/test_gatediode.sch
**.subckt test_gatediode
XM1 VD VG GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VIN VIN VG GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
VIN VIN GND dc 6.7 pulse(0 6.7 10n 10n 10n 40n 100n)
VD VD GND 1.1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/amedcalf/open-asic/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt




.option savecurrents
.control
  unset appendwrite
  save all
  op
  remzerovec
  write test_gatediode.raw
  *set appendwrite

  tran 1n 1u
  remzerovec
  write test_gatediode.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
