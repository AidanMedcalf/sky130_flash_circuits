magic
tech sky130A
magscale 1 2
timestamp 1733178670
<< error_p >>
rect -144 530 144 564
rect -174 -602 174 530
<< nwell >>
rect -144 -598 144 564
<< mvpmos >>
rect -50 -536 50 464
<< mvpdiff >>
rect -108 452 -50 464
rect -108 -524 -96 452
rect -62 -524 -50 452
rect -108 -536 -50 -524
rect 50 452 108 464
rect 50 -524 62 452
rect 96 -524 108 452
rect 50 -536 108 -524
<< mvpdiffc >>
rect -96 -524 -62 452
rect 62 -524 96 452
<< poly >>
rect -50 545 50 561
rect -50 511 -34 545
rect 34 511 50 545
rect -50 464 50 511
rect -50 -562 50 -536
<< polycont >>
rect -34 511 34 545
<< locali >>
rect -50 511 -34 545
rect 34 511 50 545
rect -96 452 -62 468
rect -96 -540 -62 -524
rect 62 452 96 468
rect 62 -540 96 -524
<< viali >>
rect -34 511 34 545
rect -96 -524 -62 452
rect 62 -524 96 452
<< metal1 >>
rect -46 545 46 551
rect -46 511 -34 545
rect 34 511 46 545
rect -46 505 46 511
rect -102 452 -56 464
rect -102 -524 -96 452
rect -62 -524 -56 452
rect -102 -536 -56 -524
rect 56 452 102 464
rect 56 -524 62 452
rect 96 -524 102 452
rect 56 -536 102 -524
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
