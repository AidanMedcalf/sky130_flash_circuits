magic
tech sky130A
magscale 1 2
timestamp 1733178670
<< error_p >>
rect -144 1030 144 1064
rect -174 -1102 174 1030
<< nwell >>
rect -144 -1098 144 1064
<< mvpmos >>
rect -50 -1036 50 964
<< mvpdiff >>
rect -108 952 -50 964
rect -108 -1024 -96 952
rect -62 -1024 -50 952
rect -108 -1036 -50 -1024
rect 50 952 108 964
rect 50 -1024 62 952
rect 96 -1024 108 952
rect 50 -1036 108 -1024
<< mvpdiffc >>
rect -96 -1024 -62 952
rect 62 -1024 96 952
<< poly >>
rect -50 1045 50 1061
rect -50 1011 -34 1045
rect 34 1011 50 1045
rect -50 964 50 1011
rect -50 -1062 50 -1036
<< polycont >>
rect -34 1011 34 1045
<< locali >>
rect -50 1011 -34 1045
rect 34 1011 50 1045
rect -96 952 -62 968
rect -96 -1040 -62 -1024
rect 62 952 96 968
rect 62 -1040 96 -1024
<< viali >>
rect -34 1011 34 1045
rect -96 -1024 -62 952
rect 62 -1024 96 952
<< metal1 >>
rect -46 1045 46 1051
rect -46 1011 -34 1045
rect 34 1011 46 1045
rect -46 1005 46 1011
rect -102 952 -56 964
rect -102 -1024 -96 952
rect -62 -1024 -56 952
rect -102 -1036 -56 -1024
rect 56 952 102 964
rect 56 -1024 62 952
rect 96 -1024 102 952
rect 56 -1036 102 -1024
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
